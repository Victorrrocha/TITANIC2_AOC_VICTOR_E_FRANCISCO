library	ieee;
use ieee.std_logic_1164.all;

entity deslocamento2bits is
	port (
	
		a 		      : in  std_logic_vector(15 downto 0);
		output      : out std_logic_vector(15 downto 0)
	);
end deslocamento2bits;

architecture implements of deslocamento2bits is 
begin 

	output <= a(13 downto 0) & "00";	
	
end implements;