LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

	entity PC is 
	port(
		A	   : in 	std_logic_vector(15 downto 0);
		Aout	: out std_logic_vector(15 downto 0)
	);
	end entity PC;

architecture adder_bh of PC is
begin 
	
	Aout <= A;
	
end adder_bh;